module top_module( output one );
    assign one = [fixme];
endmodule