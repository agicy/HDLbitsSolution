module top_module( output one );
    assign one = 1b'1;
endmodule